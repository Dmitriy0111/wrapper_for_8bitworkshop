
module example_bitmap_rom
(
    input   wire    [15 : 0]    addr, 
    output  wire    [15 : 0]    data
);
    /*******************************************************
    *               WIRE AND REG DECLARATION               *
    *******************************************************/
    reg     [15:0]      bitarray [0 : 255];
    
    assign data = bitarray[addr & 15];
    
    initial 
        $readmemb("../../fpga-examples/man.hex",bitarray);

endmodule

module sprite_scanline_renderer
#(
    parameter                   NB = 5, // 2^NB == number of sprites
    parameter                   MB = 3  // 2^MB == slots per scanline
)(
    input   wire    [0  : 0]    clk, 
    input   wire    [0  : 0]    reset, 
    input   wire    [15 : 0]    hpos, 
    input   wire    [15 : 0]    vpos, 
    output  reg     [2  : 0]    rgb,        // rgb output
    output  reg     [NB : 0]    ram_addr,   // RAM for sprite data
    input   wire    [15 : 0]    ram_data,   // (2 words per sprite)
    output  reg     [0  : 0]    ram_busy,   // set when accessing RAM
    output  reg     [15 : 0]    rom_addr,   // sprite ROM address
    input   wire    [15 : 0]    rom_data    // sprite ROM data
);
  
    localparam  N = 1 << NB, // number of sprites
                M = 1 << MB; // slots per scanline
    /*******************************************************
    *               WIRE AND REG DECLARATION               *
    *******************************************************/
    // copy of sprite data from RAM (N entries)
    reg     [7    : 0]  sprite_xpos[0 : N-1]; // X positions
    reg     [7    : 0]  sprite_ypos[0 : N-1]; // Y positions
    reg     [7    : 0]  sprite_attr[0 : N-1]; // attributes
    // M sprite slots
    reg     [7    : 0]  line_xpos[0 : M-1]; // X pos for M slots
    reg     [7    : 0]  line_yofs[0 : M-1]; // Y pos for M slots
    reg     [7    : 0]  line_attr[0 : M-1]; // attr for M slots
    reg     [0    : 0]  line_active[0 : M-1];     // slot active?
    // temporary counters
    reg     [NB-1 : 0]  i; // read index for main array (0..N-1)
    reg     [MB-1 : 0]  j; // write index for slots (0..M-1)
    reg     [MB-1 : 0]  k; // read index for slots (0..M-1)
    reg     [7    : 0]  z; // relative y offset of sprite
    reg     [8    : 0]  write_ofs; // write index of scanline buffer
    reg     [15   : 0]  out_bitmap; // shift register while writing scanline
    reg     [7    : 0]  out_attr; // attribute while writing scanline
    reg     [0    : 0]  romload; // 1 when ROM address bus is stable
    // which sprite are we currently reading?
    wire    [NB-1 : 0]  load_index;
    // RGB dual scanline buffer
    reg     [3    : 0]  scanline[0 : 511];  
    // which offset in scanline buffer to read?
    wire    [8    : 0]  read_bufidx;

    assign load_index = hpos[NB : 1];
    assign read_bufidx = { vpos[0] , hpos[7:0] };
    /*******************************************************
    *               OTHER COMB AND SEQ LOGIC               *
    *******************************************************/
    // always block (every clock cycle)
    always @(posedge clk, posedge reset)
        if( reset )
        begin
            ram_busy <= 0;
            ram_addr <= 0;
            rom_addr <= 0;
            i <= 0;
            j <= 0;
            k <= 0;
            z <= 0;
            write_ofs <= 0;
            out_bitmap <= 0;
            out_attr <= 0;
            rgb <= 0;
        end
        else
        begin
            ram_busy <= 0;
            // reset every frame, don't draw vpos >= 256
            if( vpos[8] ) 
            begin
                // load sprites from RAM on line 260
                // 8 cycles per sprite
                // do first sprite twice b/c CPU might still be busy
                if( ( vpos == 260 ) && ( hpos < N*2+8 ) ) 
                begin
                    ram_busy <= 1;
                    case( hpos[0] )
                        0: 
                        begin
                            ram_addr <= {load_index, 1'b0};
                            // load X and Y position (2 cycles ago)
                            sprite_xpos[load_index] <= ram_data[7:0];
                            sprite_ypos[load_index] <= ram_data[15:8];
                        end
                        1: 
                        begin
                            ram_addr <= {load_index, 1'b1};
                            // load attribute (2 cycles ago)
                            sprite_attr[load_index] <= ram_data[7:0];
                        end
                    endcase
                end
            end 
            else if( hpos < N*2 ) 
            begin
                // setup vars for next phase
                k <= 0;
                romload <= 0;
                // select the sprites that will appear in this scanline
                case (hpos[0])
                    // compute Y offset of sprite relative to scanline
                    0: z <= vpos - sprite_ypos[i];
                    1: begin
                        // sprite is active if Y offset is 0..15
                        if (z < 16) 
                        begin
                            line_xpos[j] <= sprite_xpos[i]; // save X pos
                            line_yofs[j] <= z; // save Y offset
                            line_attr[j] <= sprite_attr[i]; // save attr
                            line_active[j] <= 1; // mark sprite active
                            j <= j + 1; // inc counter
                        end
                        i <= i + 1; // inc main array counter
                    end
                endcase
            end 
            else if( hpos < N*2+M*18 ) 
            begin
                // setup vars for next phase
                j <= 0;
                // if sprite shift register is empty, load new sprite
                if( out_bitmap == 0 ) 
                begin
                    case( romload )
                        0: 
                        begin
                            // set ROM address and fetch bitmap
                            rom_addr <= {4'b0, line_attr[k][7:4], line_yofs[k]};
                        end
                        1: 
                        begin
                            // load scanline buffer offset to write
                            write_ofs <= {~vpos[0], line_xpos[k]};
                            // fetch 0 if sprite is inactive
                            out_bitmap <= line_active[k] ? rom_data : 0;
                            // load attribute for sprite
                            out_attr <= line_attr[k];
                            // disable sprite for next scanline
                            line_active[k] <= 0;
                            // go to next sprite in 2ndary buffer
                            k <= k + 1;
                        end
                    endcase
                    romload <= !romload;
                end else
                begin
                    // write color to scanline buffer if low bit == 1
                    if( out_bitmap[0] )
                        scanline[write_ofs] <= out_attr[3:0];
                    // shift bits right
                    out_bitmap <= out_bitmap >> 1;
                    // increment to next scanline pixel
                    write_ofs <= write_ofs + 1;
                end
            end 
            else 
            begin
                // clear counters
                i <= 0;
            end
            // read and clear buffer
            rgb <= scanline[read_bufidx];
            scanline[read_bufidx] <= 0;
        end
  
endmodule // sprite_scanline_renderer

module sprite_scanline_renderer_top
(
    input   wire    [0 : 0]     clk,
    input   wire    [0 : 0]     reset,
    output  wire    [0 : 0]     hsync,
    output  wire    [0 : 0]     vsync,
    output  wire    [2 : 0]     rgb
);
    /*******************************************************
    *                 PARAMS & LOCALPARAMS                 *
    *******************************************************/
    localparam  NB = 5,
                MB = 3;
    /*******************************************************
    *               WIRE AND REG DECLARATION               *
    *******************************************************/
    // for working with vhsync generator
    wire    [0  : 0]    display_on;         // active area
    wire    [15 : 0]    hpos;               // horizontal position from hvsync generator
    wire    [15 : 0]    vpos;               // vertical position from hvsync generator

    wire    [NB : 0]    ram_addr;
    wire    [15 : 0]    ram_data;
    wire    [0  : 0]    ram_busy;
    wire    [15 : 0]    rom_addr;
    wire    [15 : 0]    rom_data;
    wire    [2  : 0]    rgb_ssr;
    reg     [15 : 0]    ram_mem [63 : 0];
    /*******************************************************
    *                      ASSIGNMENT                      *
    *******************************************************/
    assign ram_data = ram_mem[ram_addr];
    assign rgb = { display_on,display_on,display_on } & rgb_ssr;
    /*******************************************************
    *                   MODULE INSTANCES                   *
    *******************************************************/
    // creating one hvsync generator
    hvsync_generator 
    hvsync_gen
    (
        .clk            ( clk           ),
        .reset          ( reset         ),
        .hsync          ( hsync         ),
        .vsync          ( vsync         ),
        .display_on     ( display_on    ),
        .hpos           ( hpos          ),
        .vpos           ( vpos          )
    );
    // creating one example bitmap rom
    example_bitmap_rom 
    example_bitmap_rom_0
    (
        .addr           ( rom_addr      ), 
        .data           ( rom_data      )
    );
    // creating one sprite scanline renderer
    sprite_scanline_renderer 
    #(
        .NB             ( NB            ), // 2^NB == number of sprites
        .MB             ( MB            )  // 2^MB == slots per scanline
    )
    sprite_scanline_renderer_0
    (
        .clk            ( clk           ), 
        .reset          ( reset         ), 
        .hpos           ( hpos          ), 
        .vpos           ( vpos          ), 
        .rgb            ( rgb_ssr       ),  // rgb output
        .ram_addr       ( ram_addr      ),  // RAM for sprite data
        .ram_data       ( ram_data      ),  // (2 words per sprite)
        .ram_busy       ( ram_busy      ),  // set when accessing RAM
        .rom_addr       ( rom_addr      ),  // sprite ROM address
        .rom_data       ( rom_data      )   // sprite ROM data
    );

    initial
        $readmemh( "../../fpga-examples/ram_mem.hex",ram_mem );

endmodule // sprite_scanline_renderer_top
